----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    16:22:21 02/12/2019 
-- Design Name: 
-- Module Name:    demux - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity demux is
	PORT	(
				numberA	:	IN STD_LOGIC_VECTOR(68 downto 0);
				numberB	:	IN STD_LOGIC_VECTOR(68 downto 0);
				e_data	:	IN STD_LOGIC_VECTOR(1 downto 0);
				NA0		:	OUT STD_LOGIC_VECTOR(68 downto 0);
				NB0		:	OUT STD_LOGIC_VECTOR(68 downto 0);
				NA1		:	OUT STD_LOGIC_VECTOR(68 downto 0);
				NB1		:	OUT STD_LOGIC_VECTOR(68 downto 0);
				NA2		:	OUT STD_LOGIC_VECTOR(68 downto 0);
				NB2		:	OUT STD_LOGIC_VECTOR(68 downto 0)
			);
end demux;

architecture Behavioral of demux is

begin

	PROCESS (numberA, numberB, e_data)
		begin
			case e_data is
				when "00"	=>	NA0	<=	numberA;
									NB0	<=	numberB;
									NA1	<=	"---------------------------------------------------------------------";
									NB1	<=	"---------------------------------------------------------------------";
									NA2	<=	"---------------------------------------------------------------------";
									NB2	<=	"---------------------------------------------------------------------";
				when "01"	=>	NA0	<=	"---------------------------------------------------------------------";
									NB0	<=	"---------------------------------------------------------------------";
									NA1	<=	numberA;
									NB1	<=	numberB;
									NA2	<=	"---------------------------------------------------------------------";
									NB2	<=	"---------------------------------------------------------------------";
				when "10"	=>	NA0	<=	"---------------------------------------------------------------------";
									NB0	<=	"---------------------------------------------------------------------";
									NA1	<=	"---------------------------------------------------------------------";
									NB1	<=	"---------------------------------------------------------------------";
									NA2	<=	numberA;
									NB2	<=	numberB;
				when others	=>	NA0	<=	"---------------------------------------------------------------------";
									NB0	<=	"---------------------------------------------------------------------";
									NA1	<=	"---------------------------------------------------------------------";
									NB1	<=	"---------------------------------------------------------------------";
									NA2	<=	"---------------------------------------------------------------------";
									NB2	<=	"---------------------------------------------------------------------";
				end case;
			END PROCESS;

end Behavioral;

